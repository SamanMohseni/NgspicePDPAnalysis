********************* FAP ********************
.subckt FAP VSS VDD Cout B A Cin Sum P
MMP19 Node_3 B VDD VDD PMOS
MMP4 P Node_11 Node_3 Node_3 PMOS
MMP3 Node_3 A VDD VDD PMOS
MMN19 Node_4 A VSS VSS NMOS
MMN4 P B Node_4 Node_4 NMOS
MMN3 P Node_11 VSS VSS NMOS
MMP2 Node_9 B VDD VDD PMOS
MMP1 Node_11 A Node_9 Node_9 PMOS
MMN2 Node_11 B VSS VSS NMOS
MMN1 Node_11 A VSS VSS NMOS
MMN17 Node_17 B VSS VSS NMOS
MMN16 Node_18 A Node_17 Node_17 NMOS
MMN15 Node_45 Cin Node_18 Node_18 NMOS
MMN14 Node_21 Cin VSS VSS NMOS
MMN13 Node_21 B VSS VSS NMOS
MMN12 Node_21 A VSS VSS NMOS
MMN11 Node_45 Node_19 Node_21 Node_21 NMOS
MMN9 Node_19 A Node_29 Node_29 NMOS
MMN8 Node_29 B VSS VSS NMOS
MMN7 Node_33 B VSS VSS NMOS
MMN6 Node_33 A VSS VSS NMOS
MMN5 Node_19 Cin Node_33 Node_33 NMOS
MMP9 Node_19 Cin Node_26 Node_26 PMOS
MMP8 Node_26 B VDD VDD PMOS
MMP7 Node_19 A Node_34 Node_34 PMOS
MMP6 Node_34 B Node_26 Node_26 PMOS
MMP5 Node_26 A VDD VDD PMOS
MMN10 Cout Node_19 VSS VSS NMOS
MMP10 Cout Node_19 vdd vdd PMOS
MMP11 Node_25 Cin VDD VDD PMOS
MMP12 Node_25 A VDD VDD PMOS
MMP13 Node_25 B VDD VDD PMOS
MMP14 Node_45 Node_19 Node_25 Node_25 PMOS
MMP15 Node_24 A Node_25 Node_25 PMOS
MMP16 Node_23 B Node_24 Node_24 PMOS
MMP17 Node_45 Cin Node_23 Node_23 PMOS
MMN18 Sum Node_45 VSS VSS NMOS
MMP18 Sum Node_45 VDD VDD PMOS
.ends FAP
**********************************************
